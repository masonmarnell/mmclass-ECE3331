////not used atm since I can't get the module instantiation to work right
//module DistanceSense(
//input clock,
//input LDistIn,
//input RDistIn,
//output LDistOut,
//output RDistOut

//);

////DistanceOut gets set to 1 whenever the distance sensor is triggering

////For noise suppression, a possible idea could be:
////See how many times the DistIns are giving ones withing a certain amount of clock cycles - 
//// If the count isnt high enough then don't output a 1 out of the module.

//assign LDistOut = LDistIn;
//assign RDistOut = RDistIn;

//endmodule
